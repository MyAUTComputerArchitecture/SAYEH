library IEEE;
use IEEE.std_logic_1164.all;

entity AND_COMPONENT is
	generic();
	port();
end component;

architecture AND_COMPONENT_ARCH of AND_COMPONENT is
begin

end architecture;
